//****h* rtl/common/nextCRC32_D128.vh
// NAME
//   nextCRC32_D128.vh - 
// COPYRIGHT
//   2011 - 2012 Micron Techonology, Inc.
//   Micron HMC Highly Confidential Information.
// AUTHOR
// DESCRIPTION
// HISTORY
//*****

////////////////////////////////////////////////////////////////////////////////
// Copyright (C) 1999-2008 Easics NV.
// This source file may be used and distributed without restriction
// provided that this copyright statement is not removed from the file
// and that any derivative work contains the original copyright notice
// and the associated disclaimer.
//
// THIS SOURCE FILE IS PROVIDED "AS IS" AND WITHOUT ANY EXPRESS
// OR IMPLIED WARRANTIES, INCLUDING, WITHOUT LIMITATION, THE IMPLIED
// WARRANTIES OF MERCHANTIBILITY AND FITNESS FOR A PARTICULAR PURPOSE.
//
// Purpose : synthesizable CRC function
//   * polynomial: (0 1 2 4 6 7 10 11 15 16 17 19 20 26 28 29 30 32)
//   * data width: 128
//
// Info : tools@easics.be
//        http://www.easics.com
////////////////////////////////////////////////////////////////////////////////
  function [31:0] nextCRC32_D128;

    input [127:0] Data;
    input [31:0] crc;
    reg [0:127] d;
    reg [31:0] c;
    reg [31:0] newcrc;
  begin
    d = Data;
    c = crc;

    newcrc[0] = d[126] ^ d[123] ^ d[118] ^ d[116] ^ d[115] ^ d[114] ^ d[112] ^ d[111] ^ d[108] ^ d[107] ^ d[105] ^ d[103] ^ d[102] ^ d[100] ^ d[96] ^ d[94] ^ d[92] ^ d[88] ^ d[87] ^ d[85] ^ d[83] ^ d[81] ^ d[79] ^ d[77] ^ d[75] ^ d[74] ^ d[71] ^ d[70] ^ d[68] ^ d[67] ^ d[64] ^ d[63] ^ d[62] ^ d[57] ^ d[54] ^ d[52] ^ d[51] ^ d[50] ^ d[48] ^ d[47] ^ d[46] ^ d[44] ^ d[36] ^ d[35] ^ d[34] ^ d[28] ^ d[26] ^ d[25] ^ d[24] ^ d[23] ^ d[22] ^ d[20] ^ d[17] ^ d[13] ^ d[12] ^ d[9] ^ d[7] ^ d[6] ^ d[3] ^ d[2] ^ d[0] ^ c[0] ^ c[4] ^ c[6] ^ c[7] ^ c[9] ^ c[11] ^ c[12] ^ c[15] ^ c[16] ^ c[18] ^ c[19] ^ c[20] ^ c[22] ^ c[27] ^ c[30];
    newcrc[1] = d[127] ^ d[126] ^ d[124] ^ d[123] ^ d[119] ^ d[118] ^ d[117] ^ d[114] ^ d[113] ^ d[111] ^ d[109] ^ d[107] ^ d[106] ^ d[105] ^ d[104] ^ d[102] ^ d[101] ^ d[100] ^ d[97] ^ d[96] ^ d[95] ^ d[94] ^ d[93] ^ d[92] ^ d[89] ^ d[87] ^ d[86] ^ d[85] ^ d[84] ^ d[83] ^ d[82] ^ d[81] ^ d[80] ^ d[79] ^ d[78] ^ d[77] ^ d[76] ^ d[74] ^ d[72] ^ d[70] ^ d[69] ^ d[67] ^ d[65] ^ d[62] ^ d[58] ^ d[57] ^ d[55] ^ d[54] ^ d[53] ^ d[50] ^ d[49] ^ d[46] ^ d[45] ^ d[44] ^ d[37] ^ d[34] ^ d[29] ^ d[28] ^ d[27] ^ d[22] ^ d[21] ^ d[20] ^ d[18] ^ d[17] ^ d[14] ^ d[12] ^ d[10] ^ d[9] ^ d[8] ^ d[6] ^ d[4] ^ d[2] ^ d[1] ^ d[0] ^ c[0] ^ c[1] ^ c[4] ^ c[5] ^ c[6] ^ c[8] ^ c[9] ^ c[10] ^ c[11] ^ c[13] ^ c[15] ^ c[17] ^ c[18] ^ c[21] ^ c[22] ^ c[23] ^ c[27] ^ c[28] ^ c[30] ^ c[31];
    newcrc[2] = d[127] ^ d[126] ^ d[125] ^ d[124] ^ d[123] ^ d[120] ^ d[119] ^ d[116] ^ d[111] ^ d[110] ^ d[106] ^ d[101] ^ d[100] ^ d[98] ^ d[97] ^ d[95] ^ d[93] ^ d[92] ^ d[90] ^ d[86] ^ d[84] ^ d[82] ^ d[80] ^ d[78] ^ d[74] ^ d[73] ^ d[67] ^ d[66] ^ d[64] ^ d[62] ^ d[59] ^ d[58] ^ d[57] ^ d[56] ^ d[55] ^ d[52] ^ d[48] ^ d[45] ^ d[44] ^ d[38] ^ d[36] ^ d[34] ^ d[30] ^ d[29] ^ d[26] ^ d[25] ^ d[24] ^ d[21] ^ d[20] ^ d[19] ^ d[18] ^ d[17] ^ d[15] ^ d[12] ^ d[11] ^ d[10] ^ d[6] ^ d[5] ^ d[1] ^ d[0] ^ c[1] ^ c[2] ^ c[4] ^ c[5] ^ c[10] ^ c[14] ^ c[15] ^ c[20] ^ c[23] ^ c[24] ^ c[27] ^ c[28] ^ c[29] ^ c[30] ^ c[31];
    newcrc[3] = d[127] ^ d[126] ^ d[125] ^ d[124] ^ d[121] ^ d[120] ^ d[117] ^ d[112] ^ d[111] ^ d[107] ^ d[102] ^ d[101] ^ d[99] ^ d[98] ^ d[96] ^ d[94] ^ d[93] ^ d[91] ^ d[87] ^ d[85] ^ d[83] ^ d[81] ^ d[79] ^ d[75] ^ d[74] ^ d[68] ^ d[67] ^ d[65] ^ d[63] ^ d[60] ^ d[59] ^ d[58] ^ d[57] ^ d[56] ^ d[53] ^ d[49] ^ d[46] ^ d[45] ^ d[39] ^ d[37] ^ d[35] ^ d[31] ^ d[30] ^ d[27] ^ d[26] ^ d[25] ^ d[22] ^ d[21] ^ d[20] ^ d[19] ^ d[18] ^ d[16] ^ d[13] ^ d[12] ^ d[11] ^ d[7] ^ d[6] ^ d[2] ^ d[1] ^ c[0] ^ c[2] ^ c[3] ^ c[5] ^ c[6] ^ c[11] ^ c[15] ^ c[16] ^ c[21] ^ c[24] ^ c[25] ^ c[28] ^ c[29] ^ c[30] ^ c[31];
    newcrc[4] = d[127] ^ d[125] ^ d[123] ^ d[122] ^ d[121] ^ d[116] ^ d[115] ^ d[114] ^ d[113] ^ d[111] ^ d[107] ^ d[105] ^ d[99] ^ d[97] ^ d[96] ^ d[95] ^ d[87] ^ d[86] ^ d[85] ^ d[84] ^ d[83] ^ d[82] ^ d[81] ^ d[80] ^ d[79] ^ d[77] ^ d[76] ^ d[74] ^ d[71] ^ d[70] ^ d[69] ^ d[67] ^ d[66] ^ d[63] ^ d[62] ^ d[61] ^ d[60] ^ d[59] ^ d[58] ^ d[52] ^ d[51] ^ d[48] ^ d[44] ^ d[40] ^ d[38] ^ d[35] ^ d[34] ^ d[32] ^ d[31] ^ d[27] ^ d[25] ^ d[24] ^ d[21] ^ d[19] ^ d[14] ^ d[9] ^ d[8] ^ d[6] ^ d[0] ^ c[0] ^ c[1] ^ c[3] ^ c[9] ^ c[11] ^ c[15] ^ c[17] ^ c[18] ^ c[19] ^ c[20] ^ c[25] ^ c[26] ^ c[27] ^ c[29] ^ c[31];
    newcrc[5] = d[126] ^ d[124] ^ d[123] ^ d[122] ^ d[117] ^ d[116] ^ d[115] ^ d[114] ^ d[112] ^ d[108] ^ d[106] ^ d[100] ^ d[98] ^ d[97] ^ d[96] ^ d[88] ^ d[87] ^ d[86] ^ d[85] ^ d[84] ^ d[83] ^ d[82] ^ d[81] ^ d[80] ^ d[78] ^ d[77] ^ d[75] ^ d[72] ^ d[71] ^ d[70] ^ d[68] ^ d[67] ^ d[64] ^ d[63] ^ d[62] ^ d[61] ^ d[60] ^ d[59] ^ d[53] ^ d[52] ^ d[49] ^ d[45] ^ d[41] ^ d[39] ^ d[36] ^ d[35] ^ d[33] ^ d[32] ^ d[28] ^ d[26] ^ d[25] ^ d[22] ^ d[20] ^ d[15] ^ d[10] ^ d[9] ^ d[7] ^ d[1] ^ c[0] ^ c[1] ^ c[2] ^ c[4] ^ c[10] ^ c[12] ^ c[16] ^ c[18] ^ c[19] ^ c[20] ^ c[21] ^ c[26] ^ c[27] ^ c[28] ^ c[30];
    newcrc[6] = d[127] ^ d[126] ^ d[125] ^ d[124] ^ d[117] ^ d[114] ^ d[113] ^ d[112] ^ d[111] ^ d[109] ^ d[108] ^ d[105] ^ d[103] ^ d[102] ^ d[101] ^ d[100] ^ d[99] ^ d[98] ^ d[97] ^ d[96] ^ d[94] ^ d[92] ^ d[89] ^ d[86] ^ d[84] ^ d[82] ^ d[78] ^ d[77] ^ d[76] ^ d[75] ^ d[74] ^ d[73] ^ d[72] ^ d[70] ^ d[69] ^ d[67] ^ d[65] ^ d[61] ^ d[60] ^ d[57] ^ d[53] ^ d[52] ^ d[51] ^ d[48] ^ d[47] ^ d[44] ^ d[42] ^ d[40] ^ d[37] ^ d[35] ^ d[33] ^ d[29] ^ d[28] ^ d[27] ^ d[25] ^ d[24] ^ d[22] ^ d[21] ^ d[20] ^ d[17] ^ d[16] ^ d[13] ^ d[12] ^ d[11] ^ d[10] ^ d[9] ^ d[8] ^ d[7] ^ d[6] ^ d[3] ^ d[0] ^ c[0] ^ c[1] ^ c[2] ^ c[3] ^ c[4] ^ c[5] ^ c[6] ^ c[7] ^ c[9] ^ c[12] ^ c[13] ^ c[15] ^ c[16] ^ c[17] ^ c[18] ^ c[21] ^ c[28] ^ c[29] ^ c[30] ^ c[31];
    newcrc[7] = d[127] ^ d[125] ^ d[123] ^ d[116] ^ d[113] ^ d[111] ^ d[110] ^ d[109] ^ d[108] ^ d[107] ^ d[106] ^ d[105] ^ d[104] ^ d[101] ^ d[99] ^ d[98] ^ d[97] ^ d[96] ^ d[95] ^ d[94] ^ d[93] ^ d[92] ^ d[90] ^ d[88] ^ d[81] ^ d[78] ^ d[76] ^ d[73] ^ d[67] ^ d[66] ^ d[64] ^ d[63] ^ d[61] ^ d[58] ^ d[57] ^ d[53] ^ d[51] ^ d[50] ^ d[49] ^ d[47] ^ d[46] ^ d[45] ^ d[44] ^ d[43] ^ d[41] ^ d[38] ^ d[35] ^ d[30] ^ d[29] ^ d[24] ^ d[21] ^ d[20] ^ d[18] ^ d[14] ^ d[11] ^ d[10] ^ d[8] ^ d[6] ^ d[4] ^ d[3] ^ d[2] ^ d[1] ^ d[0] ^ c[0] ^ c[1] ^ c[2] ^ c[3] ^ c[5] ^ c[8] ^ c[9] ^ c[10] ^ c[11] ^ c[12] ^ c[13] ^ c[14] ^ c[15] ^ c[17] ^ c[20] ^ c[27] ^ c[29] ^ c[31];
    newcrc[8] = d[126] ^ d[124] ^ d[117] ^ d[114] ^ d[112] ^ d[111] ^ d[110] ^ d[109] ^ d[108] ^ d[107] ^ d[106] ^ d[105] ^ d[102] ^ d[100] ^ d[99] ^ d[98] ^ d[97] ^ d[96] ^ d[95] ^ d[94] ^ d[93] ^ d[91] ^ d[89] ^ d[82] ^ d[79] ^ d[77] ^ d[74] ^ d[68] ^ d[67] ^ d[65] ^ d[64] ^ d[62] ^ d[59] ^ d[58] ^ d[54] ^ d[52] ^ d[51] ^ d[50] ^ d[48] ^ d[47] ^ d[46] ^ d[45] ^ d[44] ^ d[42] ^ d[39] ^ d[36] ^ d[31] ^ d[30] ^ d[25] ^ d[22] ^ d[21] ^ d[19] ^ d[15] ^ d[12] ^ d[11] ^ d[9] ^ d[7] ^ d[5] ^ d[4] ^ d[3] ^ d[2] ^ d[1] ^ c[0] ^ c[1] ^ c[2] ^ c[3] ^ c[4] ^ c[6] ^ c[9] ^ c[10] ^ c[11] ^ c[12] ^ c[13] ^ c[14] ^ c[15] ^ c[16] ^ c[18] ^ c[21] ^ c[28] ^ c[30];
    newcrc[9] = d[127] ^ d[125] ^ d[118] ^ d[115] ^ d[113] ^ d[112] ^ d[111] ^ d[110] ^ d[109] ^ d[108] ^ d[107] ^ d[106] ^ d[103] ^ d[101] ^ d[100] ^ d[99] ^ d[98] ^ d[97] ^ d[96] ^ d[95] ^ d[94] ^ d[92] ^ d[90] ^ d[83] ^ d[80] ^ d[78] ^ d[75] ^ d[69] ^ d[68] ^ d[66] ^ d[65] ^ d[63] ^ d[60] ^ d[59] ^ d[55] ^ d[53] ^ d[52] ^ d[51] ^ d[49] ^ d[48] ^ d[47] ^ d[46] ^ d[45] ^ d[43] ^ d[40] ^ d[37] ^ d[32] ^ d[31] ^ d[26] ^ d[23] ^ d[22] ^ d[20] ^ d[16] ^ d[13] ^ d[12] ^ d[10] ^ d[8] ^ d[6] ^ d[5] ^ d[4] ^ d[3] ^ d[2] ^ c[0] ^ c[1] ^ c[2] ^ c[3] ^ c[4] ^ c[5] ^ c[7] ^ c[10] ^ c[11] ^ c[12] ^ c[13] ^ c[14] ^ c[15] ^ c[16] ^ c[17] ^ c[19] ^ c[22] ^ c[29] ^ c[31];
    newcrc[10] = d[123] ^ d[119] ^ d[118] ^ d[115] ^ d[113] ^ d[110] ^ d[109] ^ d[105] ^ d[104] ^ d[103] ^ d[101] ^ d[99] ^ d[98] ^ d[97] ^ d[95] ^ d[94] ^ d[93] ^ d[92] ^ d[91] ^ d[88] ^ d[87] ^ d[85] ^ d[84] ^ d[83] ^ d[77] ^ d[76] ^ d[75] ^ d[74] ^ d[71] ^ d[69] ^ d[68] ^ d[66] ^ d[63] ^ d[62] ^ d[61] ^ d[60] ^ d[57] ^ d[56] ^ d[53] ^ d[51] ^ d[49] ^ d[41] ^ d[38] ^ d[36] ^ d[35] ^ d[34] ^ d[33] ^ d[32] ^ d[28] ^ d[27] ^ d[26] ^ d[25] ^ d[22] ^ d[21] ^ d[20] ^ d[14] ^ d[12] ^ d[11] ^ d[5] ^ d[4] ^ d[2] ^ d[0] ^ c[1] ^ c[2] ^ c[3] ^ c[5] ^ c[7] ^ c[8] ^ c[9] ^ c[13] ^ c[14] ^ c[17] ^ c[19] ^ c[22] ^ c[23] ^ c[27];
    newcrc[11] = d[126] ^ d[124] ^ d[123] ^ d[120] ^ d[119] ^ d[118] ^ d[115] ^ d[112] ^ d[110] ^ d[108] ^ d[107] ^ d[106] ^ d[104] ^ d[103] ^ d[99] ^ d[98] ^ d[95] ^ d[93] ^ d[89] ^ d[87] ^ d[86] ^ d[84] ^ d[83] ^ d[81] ^ d[79] ^ d[78] ^ d[76] ^ d[74] ^ d[72] ^ d[71] ^ d[69] ^ d[68] ^ d[61] ^ d[58] ^ d[51] ^ d[48] ^ d[47] ^ d[46] ^ d[44] ^ d[42] ^ d[39] ^ d[37] ^ d[33] ^ d[29] ^ d[27] ^ d[25] ^ d[24] ^ d[21] ^ d[20] ^ d[17] ^ d[15] ^ d[9] ^ d[7] ^ d[5] ^ d[2] ^ d[1] ^ d[0] ^ c[2] ^ c[3] ^ c[7] ^ c[8] ^ c[10] ^ c[11] ^ c[12] ^ c[14] ^ c[16] ^ c[19] ^ c[22] ^ c[23] ^ c[24] ^ c[27] ^ c[28] ^ c[30];
    newcrc[12] = d[127] ^ d[125] ^ d[124] ^ d[121] ^ d[120] ^ d[119] ^ d[116] ^ d[113] ^ d[111] ^ d[109] ^ d[108] ^ d[107] ^ d[105] ^ d[104] ^ d[100] ^ d[99] ^ d[96] ^ d[94] ^ d[90] ^ d[88] ^ d[87] ^ d[85] ^ d[84] ^ d[82] ^ d[80] ^ d[79] ^ d[77] ^ d[75] ^ d[73] ^ d[72] ^ d[70] ^ d[69] ^ d[62] ^ d[59] ^ d[52] ^ d[49] ^ d[48] ^ d[47] ^ d[45] ^ d[43] ^ d[40] ^ d[38] ^ d[34] ^ d[30] ^ d[28] ^ d[26] ^ d[25] ^ d[22] ^ d[21] ^ d[18] ^ d[16] ^ d[10] ^ d[8] ^ d[6] ^ d[3] ^ d[2] ^ d[1] ^ c[0] ^ c[3] ^ c[4] ^ c[8] ^ c[9] ^ c[11] ^ c[12] ^ c[13] ^ c[15] ^ c[17] ^ c[20] ^ c[23] ^ c[24] ^ c[25] ^ c[28] ^ c[29] ^ c[31];
    newcrc[13] = d[126] ^ d[125] ^ d[122] ^ d[121] ^ d[120] ^ d[117] ^ d[114] ^ d[112] ^ d[110] ^ d[109] ^ d[108] ^ d[106] ^ d[105] ^ d[101] ^ d[100] ^ d[97] ^ d[95] ^ d[91] ^ d[89] ^ d[88] ^ d[86] ^ d[85] ^ d[83] ^ d[81] ^ d[80] ^ d[78] ^ d[76] ^ d[74] ^ d[73] ^ d[71] ^ d[70] ^ d[63] ^ d[60] ^ d[53] ^ d[50] ^ d[49] ^ d[48] ^ d[46] ^ d[44] ^ d[41] ^ d[39] ^ d[35] ^ d[31] ^ d[29] ^ d[27] ^ d[26] ^ d[23] ^ d[22] ^ d[19] ^ d[17] ^ d[11] ^ d[9] ^ d[7] ^ d[4] ^ d[3] ^ d[2] ^ c[1] ^ c[4] ^ c[5] ^ c[9] ^ c[10] ^ c[12] ^ c[13] ^ c[14] ^ c[16] ^ c[18] ^ c[21] ^ c[24] ^ c[25] ^ c[26] ^ c[29] ^ c[30];
    newcrc[14] = d[127] ^ d[126] ^ d[123] ^ d[122] ^ d[121] ^ d[118] ^ d[115] ^ d[113] ^ d[111] ^ d[110] ^ d[109] ^ d[107] ^ d[106] ^ d[102] ^ d[101] ^ d[98] ^ d[96] ^ d[92] ^ d[90] ^ d[89] ^ d[87] ^ d[86] ^ d[84] ^ d[82] ^ d[81] ^ d[79] ^ d[77] ^ d[75] ^ d[74] ^ d[72] ^ d[71] ^ d[64] ^ d[61] ^ d[54] ^ d[51] ^ d[50] ^ d[49] ^ d[47] ^ d[45] ^ d[42] ^ d[40] ^ d[36] ^ d[32] ^ d[30] ^ d[28] ^ d[27] ^ d[24] ^ d[23] ^ d[20] ^ d[18] ^ d[12] ^ d[10] ^ d[8] ^ d[5] ^ d[4] ^ d[3] ^ c[0] ^ c[2] ^ c[5] ^ c[6] ^ c[10] ^ c[11] ^ c[13] ^ c[14] ^ c[15] ^ c[17] ^ c[19] ^ c[22] ^ c[25] ^ c[26] ^ c[27] ^ c[30] ^ c[31];
    newcrc[15] = d[127] ^ d[126] ^ d[124] ^ d[122] ^ d[119] ^ d[118] ^ d[115] ^ d[110] ^ d[105] ^ d[100] ^ d[99] ^ d[97] ^ d[96] ^ d[94] ^ d[93] ^ d[92] ^ d[91] ^ d[90] ^ d[82] ^ d[81] ^ d[80] ^ d[79] ^ d[78] ^ d[77] ^ d[76] ^ d[74] ^ d[73] ^ d[72] ^ d[71] ^ d[70] ^ d[68] ^ d[67] ^ d[65] ^ d[64] ^ d[63] ^ d[57] ^ d[55] ^ d[54] ^ d[47] ^ d[44] ^ d[43] ^ d[41] ^ d[37] ^ d[36] ^ d[35] ^ d[34] ^ d[33] ^ d[31] ^ d[29] ^ d[26] ^ d[23] ^ d[22] ^ d[21] ^ d[20] ^ d[19] ^ d[17] ^ d[12] ^ d[11] ^ d[7] ^ d[5] ^ d[4] ^ d[3] ^ d[2] ^ d[0] ^ c[0] ^ c[1] ^ c[3] ^ c[4] ^ c[9] ^ c[14] ^ c[19] ^ c[22] ^ c[23] ^ c[26] ^ c[28] ^ c[30] ^ c[31];
    newcrc[16] = d[127] ^ d[126] ^ d[125] ^ d[120] ^ d[119] ^ d[118] ^ d[115] ^ d[114] ^ d[112] ^ d[108] ^ d[107] ^ d[106] ^ d[105] ^ d[103] ^ d[102] ^ d[101] ^ d[98] ^ d[97] ^ d[96] ^ d[95] ^ d[93] ^ d[91] ^ d[88] ^ d[87] ^ d[85] ^ d[82] ^ d[80] ^ d[78] ^ d[73] ^ d[72] ^ d[70] ^ d[69] ^ d[67] ^ d[66] ^ d[65] ^ d[63] ^ d[62] ^ d[58] ^ d[57] ^ d[56] ^ d[55] ^ d[54] ^ d[52] ^ d[51] ^ d[50] ^ d[47] ^ d[46] ^ d[45] ^ d[42] ^ d[38] ^ d[37] ^ d[32] ^ d[30] ^ d[28] ^ d[27] ^ d[26] ^ d[25] ^ d[21] ^ d[18] ^ d[17] ^ d[9] ^ d[8] ^ d[7] ^ d[5] ^ d[4] ^ d[2] ^ d[1] ^ d[0] ^ c[0] ^ c[1] ^ c[2] ^ c[5] ^ c[6] ^ c[7] ^ c[9] ^ c[10] ^ c[11] ^ c[12] ^ c[16] ^ c[18] ^ c[19] ^ c[22] ^ c[23] ^ c[24] ^ c[29] ^ c[30] ^ c[31];
    newcrc[17] = d[127] ^ d[123] ^ d[121] ^ d[120] ^ d[119] ^ d[118] ^ d[114] ^ d[113] ^ d[112] ^ d[111] ^ d[109] ^ d[106] ^ d[105] ^ d[104] ^ d[100] ^ d[99] ^ d[98] ^ d[97] ^ d[89] ^ d[87] ^ d[86] ^ d[85] ^ d[77] ^ d[75] ^ d[73] ^ d[66] ^ d[62] ^ d[59] ^ d[58] ^ d[56] ^ d[55] ^ d[54] ^ d[53] ^ d[50] ^ d[44] ^ d[43] ^ d[39] ^ d[38] ^ d[36] ^ d[35] ^ d[34] ^ d[33] ^ d[31] ^ d[29] ^ d[27] ^ d[25] ^ d[24] ^ d[23] ^ d[20] ^ d[19] ^ d[18] ^ d[17] ^ d[13] ^ d[12] ^ d[10] ^ d[8] ^ d[7] ^ d[5] ^ d[1] ^ d[0] ^ c[1] ^ c[2] ^ c[3] ^ c[4] ^ c[8] ^ c[9] ^ c[10] ^ c[13] ^ c[15] ^ c[16] ^ c[17] ^ c[18] ^ c[22] ^ c[23] ^ c[24] ^ c[25] ^ c[27] ^ c[31];
    newcrc[18] = d[124] ^ d[122] ^ d[121] ^ d[120] ^ d[119] ^ d[115] ^ d[114] ^ d[113] ^ d[112] ^ d[110] ^ d[107] ^ d[106] ^ d[105] ^ d[101] ^ d[100] ^ d[99] ^ d[98] ^ d[90] ^ d[88] ^ d[87] ^ d[86] ^ d[78] ^ d[76] ^ d[74] ^ d[67] ^ d[63] ^ d[60] ^ d[59] ^ d[57] ^ d[56] ^ d[55] ^ d[54] ^ d[51] ^ d[45] ^ d[44] ^ d[40] ^ d[39] ^ d[37] ^ d[36] ^ d[35] ^ d[34] ^ d[32] ^ d[30] ^ d[28] ^ d[26] ^ d[25] ^ d[24] ^ d[21] ^ d[20] ^ d[19] ^ d[18] ^ d[14] ^ d[13] ^ d[11] ^ d[9] ^ d[8] ^ d[6] ^ d[2] ^ d[1] ^ c[2] ^ c[3] ^ c[4] ^ c[5] ^ c[9] ^ c[10] ^ c[11] ^ c[14] ^ c[16] ^ c[17] ^ c[18] ^ c[19] ^ c[23] ^ c[24] ^ c[25] ^ c[26] ^ c[28];
    newcrc[19] = d[126] ^ d[125] ^ d[122] ^ d[121] ^ d[120] ^ d[118] ^ d[113] ^ d[112] ^ d[106] ^ d[105] ^ d[103] ^ d[101] ^ d[99] ^ d[96] ^ d[94] ^ d[92] ^ d[91] ^ d[89] ^ d[85] ^ d[83] ^ d[81] ^ d[74] ^ d[71] ^ d[70] ^ d[67] ^ d[63] ^ d[62] ^ d[61] ^ d[60] ^ d[58] ^ d[56] ^ d[55] ^ d[54] ^ d[51] ^ d[50] ^ d[48] ^ d[47] ^ d[45] ^ d[44] ^ d[41] ^ d[40] ^ d[38] ^ d[37] ^ d[34] ^ d[33] ^ d[31] ^ d[29] ^ d[28] ^ d[27] ^ d[24] ^ d[23] ^ d[21] ^ d[19] ^ d[17] ^ d[15] ^ d[14] ^ d[13] ^ d[10] ^ d[6] ^ d[0] ^ c[0] ^ c[3] ^ c[5] ^ c[7] ^ c[9] ^ c[10] ^ c[16] ^ c[17] ^ c[22] ^ c[24] ^ c[25] ^ c[26] ^ c[29] ^ c[30];
    newcrc[20] = d[127] ^ d[122] ^ d[121] ^ d[119] ^ d[118] ^ d[116] ^ d[115] ^ d[113] ^ d[112] ^ d[111] ^ d[108] ^ d[106] ^ d[105] ^ d[104] ^ d[103] ^ d[97] ^ d[96] ^ d[95] ^ d[94] ^ d[93] ^ d[90] ^ d[88] ^ d[87] ^ d[86] ^ d[85] ^ d[84] ^ d[83] ^ d[82] ^ d[81] ^ d[79] ^ d[77] ^ d[74] ^ d[72] ^ d[70] ^ d[67] ^ d[61] ^ d[59] ^ d[56] ^ d[55] ^ d[54] ^ d[50] ^ d[49] ^ d[47] ^ d[45] ^ d[44] ^ d[42] ^ d[41] ^ d[39] ^ d[38] ^ d[36] ^ d[32] ^ d[30] ^ d[29] ^ d[26] ^ d[23] ^ d[18] ^ d[17] ^ d[16] ^ d[15] ^ d[14] ^ d[13] ^ d[12] ^ d[11] ^ d[9] ^ d[6] ^ d[3] ^ d[2] ^ d[1] ^ d[0] ^ c[0] ^ c[1] ^ c[7] ^ c[8] ^ c[9] ^ c[10] ^ c[12] ^ c[15] ^ c[16] ^ c[17] ^ c[19] ^ c[20] ^ c[22] ^ c[23] ^ c[25] ^ c[26] ^ c[31];
    newcrc[21] = d[123] ^ d[122] ^ d[120] ^ d[119] ^ d[117] ^ d[116] ^ d[114] ^ d[113] ^ d[112] ^ d[109] ^ d[107] ^ d[106] ^ d[105] ^ d[104] ^ d[98] ^ d[97] ^ d[96] ^ d[95] ^ d[94] ^ d[91] ^ d[89] ^ d[88] ^ d[87] ^ d[86] ^ d[85] ^ d[84] ^ d[83] ^ d[82] ^ d[80] ^ d[78] ^ d[75] ^ d[73] ^ d[71] ^ d[68] ^ d[62] ^ d[60] ^ d[57] ^ d[56] ^ d[55] ^ d[51] ^ d[50] ^ d[48] ^ d[46] ^ d[45] ^ d[43] ^ d[42] ^ d[40] ^ d[39] ^ d[37] ^ d[33] ^ d[31] ^ d[30] ^ d[27] ^ d[24] ^ d[19] ^ d[18] ^ d[17] ^ d[16] ^ d[15] ^ d[14] ^ d[13] ^ d[12] ^ d[10] ^ d[7] ^ d[4] ^ d[3] ^ d[2] ^ d[1] ^ c[0] ^ c[1] ^ c[2] ^ c[8] ^ c[9] ^ c[10] ^ c[11] ^ c[13] ^ c[16] ^ c[17] ^ c[18] ^ c[20] ^ c[21] ^ c[23] ^ c[24] ^ c[26] ^ c[27];
    newcrc[22] = d[124] ^ d[123] ^ d[121] ^ d[120] ^ d[118] ^ d[117] ^ d[115] ^ d[114] ^ d[113] ^ d[110] ^ d[108] ^ d[107] ^ d[106] ^ d[105] ^ d[99] ^ d[98] ^ d[97] ^ d[96] ^ d[95] ^ d[92] ^ d[90] ^ d[89] ^ d[88] ^ d[87] ^ d[86] ^ d[85] ^ d[84] ^ d[83] ^ d[81] ^ d[79] ^ d[76] ^ d[74] ^ d[72] ^ d[69] ^ d[63] ^ d[61] ^ d[58] ^ d[57] ^ d[56] ^ d[52] ^ d[51] ^ d[49] ^ d[47] ^ d[46] ^ d[44] ^ d[43] ^ d[41] ^ d[40] ^ d[38] ^ d[34] ^ d[32] ^ d[31] ^ d[28] ^ d[25] ^ d[20] ^ d[19] ^ d[18] ^ d[17] ^ d[16] ^ d[15] ^ d[14] ^ d[13] ^ d[11] ^ d[8] ^ d[5] ^ d[4] ^ d[3] ^ d[2] ^ c[0] ^ c[1] ^ c[2] ^ c[3] ^ c[9] ^ c[10] ^ c[11] ^ c[12] ^ c[14] ^ c[17] ^ c[18] ^ c[19] ^ c[21] ^ c[22] ^ c[24] ^ c[25] ^ c[27] ^ c[28];
    newcrc[23] = d[125] ^ d[124] ^ d[122] ^ d[121] ^ d[119] ^ d[118] ^ d[116] ^ d[115] ^ d[114] ^ d[111] ^ d[109] ^ d[108] ^ d[107] ^ d[106] ^ d[100] ^ d[99] ^ d[98] ^ d[97] ^ d[96] ^ d[93] ^ d[91] ^ d[90] ^ d[89] ^ d[88] ^ d[87] ^ d[86] ^ d[85] ^ d[84] ^ d[82] ^ d[80] ^ d[77] ^ d[75] ^ d[73] ^ d[70] ^ d[64] ^ d[62] ^ d[59] ^ d[58] ^ d[57] ^ d[53] ^ d[52] ^ d[50] ^ d[48] ^ d[47] ^ d[45] ^ d[44] ^ d[42] ^ d[41] ^ d[39] ^ d[35] ^ d[33] ^ d[32] ^ d[29] ^ d[26] ^ d[21] ^ d[20] ^ d[19] ^ d[18] ^ d[17] ^ d[16] ^ d[15] ^ d[14] ^ d[12] ^ d[9] ^ d[6] ^ d[5] ^ d[4] ^ d[3] ^ c[0] ^ c[1] ^ c[2] ^ c[3] ^ c[4] ^ c[10] ^ c[11] ^ c[12] ^ c[13] ^ c[15] ^ c[18] ^ c[19] ^ c[20] ^ c[22] ^ c[23] ^ c[25] ^ c[26] ^ c[28] ^ c[29];
    newcrc[24] = d[126] ^ d[125] ^ d[123] ^ d[122] ^ d[120] ^ d[119] ^ d[117] ^ d[116] ^ d[115] ^ d[112] ^ d[110] ^ d[109] ^ d[108] ^ d[107] ^ d[101] ^ d[100] ^ d[99] ^ d[98] ^ d[97] ^ d[94] ^ d[92] ^ d[91] ^ d[90] ^ d[89] ^ d[88] ^ d[87] ^ d[86] ^ d[85] ^ d[83] ^ d[81] ^ d[78] ^ d[76] ^ d[74] ^ d[71] ^ d[65] ^ d[63] ^ d[60] ^ d[59] ^ d[58] ^ d[54] ^ d[53] ^ d[51] ^ d[49] ^ d[48] ^ d[46] ^ d[45] ^ d[43] ^ d[42] ^ d[40] ^ d[36] ^ d[34] ^ d[33] ^ d[30] ^ d[27] ^ d[22] ^ d[21] ^ d[20] ^ d[19] ^ d[18] ^ d[17] ^ d[16] ^ d[15] ^ d[13] ^ d[10] ^ d[7] ^ d[6] ^ d[5] ^ d[4] ^ c[1] ^ c[2] ^ c[3] ^ c[4] ^ c[5] ^ c[11] ^ c[12] ^ c[13] ^ c[14] ^ c[16] ^ c[19] ^ c[20] ^ c[21] ^ c[23] ^ c[24] ^ c[26] ^ c[27] ^ c[29] ^ c[30];
    newcrc[25] = d[127] ^ d[126] ^ d[124] ^ d[123] ^ d[121] ^ d[120] ^ d[118] ^ d[117] ^ d[116] ^ d[113] ^ d[111] ^ d[110] ^ d[109] ^ d[108] ^ d[102] ^ d[101] ^ d[100] ^ d[99] ^ d[98] ^ d[95] ^ d[93] ^ d[92] ^ d[91] ^ d[90] ^ d[89] ^ d[88] ^ d[87] ^ d[86] ^ d[84] ^ d[82] ^ d[79] ^ d[77] ^ d[75] ^ d[72] ^ d[66] ^ d[64] ^ d[61] ^ d[60] ^ d[59] ^ d[55] ^ d[54] ^ d[52] ^ d[50] ^ d[49] ^ d[47] ^ d[46] ^ d[44] ^ d[43] ^ d[41] ^ d[37] ^ d[35] ^ d[34] ^ d[31] ^ d[28] ^ d[23] ^ d[22] ^ d[21] ^ d[20] ^ d[19] ^ d[18] ^ d[17] ^ d[16] ^ d[14] ^ d[11] ^ d[8] ^ d[7] ^ d[6] ^ d[5] ^ c[2] ^ c[3] ^ c[4] ^ c[5] ^ c[6] ^ c[12] ^ c[13] ^ c[14] ^ c[15] ^ c[17] ^ c[20] ^ c[21] ^ c[22] ^ c[24] ^ c[25] ^ c[27] ^ c[28] ^ c[30] ^ c[31];
    newcrc[26] = d[127] ^ d[126] ^ d[125] ^ d[124] ^ d[123] ^ d[122] ^ d[121] ^ d[119] ^ d[117] ^ d[116] ^ d[115] ^ d[110] ^ d[109] ^ d[108] ^ d[107] ^ d[105] ^ d[101] ^ d[99] ^ d[93] ^ d[91] ^ d[90] ^ d[89] ^ d[81] ^ d[80] ^ d[79] ^ d[78] ^ d[77] ^ d[76] ^ d[75] ^ d[74] ^ d[73] ^ d[71] ^ d[70] ^ d[68] ^ d[65] ^ d[64] ^ d[63] ^ d[61] ^ d[60] ^ d[57] ^ d[56] ^ d[55] ^ d[54] ^ d[53] ^ d[52] ^ d[46] ^ d[45] ^ d[42] ^ d[38] ^ d[34] ^ d[32] ^ d[29] ^ d[28] ^ d[26] ^ d[25] ^ d[21] ^ d[19] ^ d[18] ^ d[15] ^ d[13] ^ d[8] ^ d[3] ^ d[2] ^ d[0] ^ c[3] ^ c[5] ^ c[9] ^ c[11] ^ c[12] ^ c[13] ^ c[14] ^ c[19] ^ c[20] ^ c[21] ^ c[23] ^ c[25] ^ c[26] ^ c[27] ^ c[28] ^ c[29] ^ c[30] ^ c[31];
    newcrc[27] = d[127] ^ d[126] ^ d[125] ^ d[124] ^ d[123] ^ d[122] ^ d[120] ^ d[118] ^ d[117] ^ d[116] ^ d[111] ^ d[110] ^ d[109] ^ d[108] ^ d[106] ^ d[102] ^ d[100] ^ d[94] ^ d[92] ^ d[91] ^ d[90] ^ d[82] ^ d[81] ^ d[80] ^ d[79] ^ d[78] ^ d[77] ^ d[76] ^ d[75] ^ d[74] ^ d[72] ^ d[71] ^ d[69] ^ d[66] ^ d[65] ^ d[64] ^ d[62] ^ d[61] ^ d[58] ^ d[57] ^ d[56] ^ d[55] ^ d[54] ^ d[53] ^ d[47] ^ d[46] ^ d[43] ^ d[39] ^ d[35] ^ d[33] ^ d[30] ^ d[29] ^ d[27] ^ d[26] ^ d[22] ^ d[20] ^ d[19] ^ d[16] ^ d[14] ^ d[9] ^ d[4] ^ d[3] ^ d[1] ^ c[4] ^ c[6] ^ c[10] ^ c[12] ^ c[13] ^ c[14] ^ c[15] ^ c[20] ^ c[21] ^ c[22] ^ c[24] ^ c[26] ^ c[27] ^ c[28] ^ c[29] ^ c[30] ^ c[31];
    newcrc[28] = d[127] ^ d[125] ^ d[124] ^ d[121] ^ d[119] ^ d[117] ^ d[116] ^ d[115] ^ d[114] ^ d[110] ^ d[109] ^ d[108] ^ d[105] ^ d[102] ^ d[101] ^ d[100] ^ d[96] ^ d[95] ^ d[94] ^ d[93] ^ d[91] ^ d[88] ^ d[87] ^ d[85] ^ d[82] ^ d[80] ^ d[78] ^ d[76] ^ d[74] ^ d[73] ^ d[72] ^ d[71] ^ d[68] ^ d[66] ^ d[65] ^ d[64] ^ d[59] ^ d[58] ^ d[56] ^ d[55] ^ d[52] ^ d[51] ^ d[50] ^ d[46] ^ d[40] ^ d[35] ^ d[31] ^ d[30] ^ d[27] ^ d[26] ^ d[25] ^ d[24] ^ d[22] ^ d[21] ^ d[15] ^ d[13] ^ d[12] ^ d[10] ^ d[9] ^ d[7] ^ d[6] ^ d[5] ^ d[4] ^ d[3] ^ d[0] ^ c[0] ^ c[4] ^ c[5] ^ c[6] ^ c[9] ^ c[12] ^ c[13] ^ c[14] ^ c[18] ^ c[19] ^ c[20] ^ c[21] ^ c[23] ^ c[25] ^ c[28] ^ c[29] ^ c[31];
    newcrc[29] = d[125] ^ d[123] ^ d[122] ^ d[120] ^ d[117] ^ d[114] ^ d[112] ^ d[110] ^ d[109] ^ d[108] ^ d[107] ^ d[106] ^ d[105] ^ d[101] ^ d[100] ^ d[97] ^ d[95] ^ d[89] ^ d[87] ^ d[86] ^ d[85] ^ d[73] ^ d[72] ^ d[71] ^ d[70] ^ d[69] ^ d[68] ^ d[66] ^ d[65] ^ d[64] ^ d[63] ^ d[62] ^ d[60] ^ d[59] ^ d[56] ^ d[54] ^ d[53] ^ d[50] ^ d[48] ^ d[46] ^ d[44] ^ d[41] ^ d[35] ^ d[34] ^ d[32] ^ d[31] ^ d[27] ^ d[24] ^ d[20] ^ d[17] ^ d[16] ^ d[14] ^ d[12] ^ d[11] ^ d[10] ^ d[9] ^ d[8] ^ d[5] ^ d[4] ^ d[3] ^ d[2] ^ d[1] ^ d[0] ^ c[1] ^ c[4] ^ c[5] ^ c[9] ^ c[10] ^ c[11] ^ c[12] ^ c[13] ^ c[14] ^ c[16] ^ c[18] ^ c[21] ^ c[24] ^ c[26] ^ c[27] ^ c[29];
    newcrc[30] = d[124] ^ d[121] ^ d[116] ^ d[114] ^ d[113] ^ d[112] ^ d[110] ^ d[109] ^ d[106] ^ d[105] ^ d[103] ^ d[101] ^ d[100] ^ d[98] ^ d[94] ^ d[92] ^ d[90] ^ d[86] ^ d[85] ^ d[83] ^ d[81] ^ d[79] ^ d[77] ^ d[75] ^ d[73] ^ d[72] ^ d[69] ^ d[68] ^ d[66] ^ d[65] ^ d[62] ^ d[61] ^ d[60] ^ d[55] ^ d[52] ^ d[50] ^ d[49] ^ d[48] ^ d[46] ^ d[45] ^ d[44] ^ d[42] ^ d[34] ^ d[33] ^ d[32] ^ d[26] ^ d[24] ^ d[23] ^ d[22] ^ d[21] ^ d[20] ^ d[18] ^ d[15] ^ d[11] ^ d[10] ^ d[7] ^ d[5] ^ d[4] ^ d[1] ^ d[0] ^ c[2] ^ c[4] ^ c[5] ^ c[7] ^ c[9] ^ c[10] ^ c[13] ^ c[14] ^ c[16] ^ c[17] ^ c[18] ^ c[20] ^ c[25] ^ c[28];
    newcrc[31] = d[125] ^ d[122] ^ d[117] ^ d[115] ^ d[114] ^ d[113] ^ d[111] ^ d[110] ^ d[107] ^ d[106] ^ d[104] ^ d[102] ^ d[101] ^ d[99] ^ d[95] ^ d[93] ^ d[91] ^ d[87] ^ d[86] ^ d[84] ^ d[82] ^ d[80] ^ d[78] ^ d[76] ^ d[74] ^ d[73] ^ d[70] ^ d[69] ^ d[67] ^ d[66] ^ d[63] ^ d[62] ^ d[61] ^ d[56] ^ d[53] ^ d[51] ^ d[50] ^ d[49] ^ d[47] ^ d[46] ^ d[45] ^ d[43] ^ d[35] ^ d[34] ^ d[33] ^ d[27] ^ d[25] ^ d[24] ^ d[23] ^ d[22] ^ d[21] ^ d[19] ^ d[16] ^ d[12] ^ d[11] ^ d[8] ^ d[6] ^ d[5] ^ d[2] ^ d[1] ^ c[3] ^ c[5] ^ c[6] ^ c[8] ^ c[10] ^ c[11] ^ c[14] ^ c[15] ^ c[17] ^ c[18] ^ c[19] ^ c[21] ^ c[26] ^ c[29];
    nextCRC32_D128 = newcrc;
  end
  endfunction
